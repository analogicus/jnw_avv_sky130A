*Automatic generated instance fron ../../tech/scripts/gensvinst tmpDig
adut [clk
+ reset
+ cmp
+ tmpPulse
+ ]
+ [PI1
+ PI2
+ PII1
+ dummy
+ PII2
+ PA
+ PB
+ PC
+ PD
+ s_BG2CMP
+ s_BgCtrl
+ s_PtatCtrl
+ s_Cap2CMP
+ s_Ref2CMP
+ s_CapRst
+ s_PtatOut
+ s_Rdiscon_N
+ s_CmpOutDisable
+ src_n
+ snk
+ cmp_p1
+ cmp_p2
+ PwrUp
+ rst
+ valid
+ preChrg
+ setupBias
+ tmpCount_out.7
+ tmpCount_out.6
+ tmpCount_out.5
+ tmpCount_out.4
+ tmpCount_out.3
+ tmpCount_out.2
+ tmpCount_out.1
+ tmpCount_out.0
+ ] null dut
.model dut d_cosim simulation="../tmpDig.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 reset 0 1G
Rsvi2 cmp 0 1G
Rsvi3 tmpPulse 0 1G

* Outputs
Rsvi4 PI1 0 1G
Rsvi5 PI2 0 1G
Rsvi6 PII1 0 1G
Rsvi7 dummy 0 1G
Rsvi8 PII2 0 1G
Rsvi9 PA 0 1G
Rsvi10 PB 0 1G
Rsvi11 PC 0 1G
Rsvi12 PD 0 1G
Rsvi13 s_BG2CMP 0 1G
Rsvi14 s_BgCtrl 0 1G
Rsvi15 s_PtatCtrl 0 1G
Rsvi16 s_Cap2CMP 0 1G
Rsvi17 s_Ref2CMP 0 1G
Rsvi18 s_CapRst 0 1G
Rsvi19 s_PtatOut 0 1G
Rsvi20 s_Rdiscon_N 0 1G
Rsvi21 s_CmpOutDisable 0 1G
Rsvi22 src_n 0 1G
Rsvi23 snk 0 1G
Rsvi24 cmp_p1 0 1G
Rsvi25 cmp_p2 0 1G
Rsvi26 PwrUp 0 1G
Rsvi27 rst 0 1G
Rsvi28 valid 0 1G
Rsvi29 preChrg 0 1G
Rsvi30 setupBias 0 1G
Rsvi31 tmpCount_out.7 0 1G
Rsvi32 tmpCount_out.6 0 1G
Rsvi33 tmpCount_out.5 0 1G
Rsvi34 tmpCount_out.4 0 1G
Rsvi35 tmpCount_out.3 0 1G
Rsvi36 tmpCount_out.2 0 1G
Rsvi37 tmpCount_out.1 0 1G
Rsvi38 tmpCount_out.0 0 1G

.save v(PI1)

.save v(PI2)

.save v(PII1)

.save v(dummy)

.save v(PII2)

.save v(PA)

.save v(PB)

.save v(PC)

.save v(PD)

.save v(s_BG2CMP)

.save v(s_BgCtrl)

.save v(s_PtatCtrl)

.save v(s_Cap2CMP)

.save v(s_Ref2CMP)

.save v(s_CapRst)

.save v(s_PtatOut)

.save v(s_Rdiscon_N)

.save v(s_CmpOutDisable)

.save v(src_n)

.save v(snk)

.save v(cmp_p1)

.save v(cmp_p2)

.save v(PwrUp)

.save v(rst)

.save v(valid)

.save v(preChrg)

.save v(setupBias)

E_STATE_tmpCount_out dec_tmpCount_out 0 value={( 0 
+ + 128*v(tmpCount_out.7)/AVDD
+ + 64*v(tmpCount_out.6)/AVDD
+ + 32*v(tmpCount_out.5)/AVDD
+ + 16*v(tmpCount_out.4)/AVDD
+ + 8*v(tmpCount_out.3)/AVDD
+ + 4*v(tmpCount_out.2)/AVDD
+ + 2*v(tmpCount_out.1)/AVDD
+ + 1*v(tmpCount_out.0)/AVDD
+)/1000}
.save v(dec_tmpCount_out)

