*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bgTest_lpe.spi
#else
.include ../../../work/xsch/bgTest.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=25 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc 1.8

* VA  A  0  pulse(0 1.8 0 10p 10p 50n 100n)
VB  B  0  pulse(0.8 1.1 0 10p 10p 100n 200n)
* VA  A  0  pwl 0 0 50n 0 51n 1.8 150n 1.8 151n 0
* VB  B  0  pwl 0 0 100n 0 101n 1.8 200n 1.8 201n 0




*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(vdd)
.save v(vss)
.save i(xdut.v_itot)
.save i(xdut.v_ip1)
.save i(xdut.v_ip2)
.save i(xdut.v_in1)
.save i(xdut.v_in2)
.save v(vref)
.save v(vp)
.save v(vn)
.save v(xdut.vctrl)
.save v(VBE)
.save v(A)
.save v(B)
.save v(xdut.y)
.save v(xdut.clk1)
.save v(xdut.clk2)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


*dc TEMP -40 125 1
set fend = .raw


* foreach vtemp -40 40 120
*   option temp=$vtemp
*   tran 1n 500n
*   write {cicname}_$vtemp$fend
* end

tran 1n 500n

write
quit


.endc

.end
