*cicsimgen tran

.param SEED=0

*Nothing here

.param mc_mm_switch=0
.param mc_pr_switch=0
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__ss.pm3.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__ss.corner.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.tech/ngspice/corners/ss/nonfet.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.tech/ngspice/all.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.tech/ngspice/r+c/res_high__cap_high.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.tech/ngspice/r+c/res_high__cap_high__lin.spice"
.include "/cad/gnu/oseda/sky130nm/2024-08/share/pdk/sky130A/libs.tech/ngspice/corners/ss/specialized_cells.spice"

.lib "../../../tech/ngspice/temperature.spi" Tt

.lib "../../../tech/ngspice/supply.spi" Vh

*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../work/xsch/TB_bandgap.spice



*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option GMIN=1e-15 TNOM=25 
* .option TEMP=25

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {1.8}
.param PERIOD_CLK = {50e-9}
.param PW_CLK = PERIOD_CLK/2
.param T_START = PERIOD_CLK*4
.param T_RESET = {T_START + PERIOD_CLK + PW_CLK}
.param T_RESET_F = {T_RESET + 1n}
.param nbpt = 9*(8+5+2)

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS    0   dc 0
VDD  vdd    0   dc 1.8
VRST reset  0   dc 0
VCLK clk    0   dc 0 pulse (0 {AVDD} {T_START} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(clk)
.save v(vdd)
.save v(vss)
.save v(pa)
.save v(pb)
.save v(pc)
.save v(pd)
.save v(pi1)
.save v(pi2)
.save v(pii1)
.save v(pii2)
.save v(vref)
.save v(valid)
.save v(snk)
.save v(src)
.save v(xdut.vctrl)
.save v(xdut.pbias)
.save v(xdut.nbias)
.save v(xdut.vp)
.save v(xdut.vn)
.save v(reset)
.save v(rst)
.save v(cmp)
.save v(xdut.x3.snk_gate)
.save v(xdut.x3.src_gate_n)
.save v(xdut.x3.src_cap)
.save v(xdut.x3.snk_cap)
.save i(xdut.v_nbias)
.save i(xdut.v_pbias)
.save i(xdut.x2.vipmos)
.save v(xdut.x2.Hcharge)
.save v(xdut.x2.Lcharge)
.save v(xdut.x2.outRes)
.save v(xdut.x3.Vpre)


* .save all
* .option savecurrents


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

unset askquit

optran 0 0 0 100p 1.5u 0


set fend = .raw


* tran 70n 40u

foreach vtemp -40 20 80 125
  option temp=$vtemp
  tran 1000n 60u
  write tran_SchGtKssTtVh_$vtemp$fend
end

* foreach vtemp -40 -39 -38 -37 -36 -34 -32 -30 -28 -26 -24 -22 -20 -18 -16 -14 -12 -10 -8 -6 -4 -2 0 20 40 50
*   .save all
*   option temp=$vtemp
*   option savecurrents
*   tran 1000n 80u
*   write tran_SchGtKssTtVh_debug_$vtemp$fend
* end


write
quit


.endc

.end

