*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_charge_pump_lpe.spi
#else
.include ../../../work/xsch/TB_charge_pump.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=20 GMIN=1e-15

.param TRF = 10p
.param AVDD = {1.8}
.param PERIOD_CLK = {50e-9}
.param PW_CLK = PERIOD_CLK/2
.param T_START = PERIOD_CLK*4
.param T_RESET = {T_START + PERIOD_CLK + PW_CLK}
.param T_RESET_F = {T_RESET + 1n}
.param nbpt = 9*(8+5+2)

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS    0   dc 0
VDD  vdd    0   dc 1.8
VRST reset  0   dc 0
VCLK clk    0   dc 0 pulse (0 {AVDD} {T_START} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(vdd) 
.save v(vss)
.save v(src_n)
.save v(snk)
.save v(vctrl)
.save v(xdut.pbias)
.save v(xdut.nbias)
.save v(preChrg)
.save v(xdut.x1.snk_gate)
.save v(xdut.x1.src_gate_n)
.save v(xdut.x1.src_cap)
.save v(xdut.x1.snk_cap)
.save i(xdut.x1.v_isrc)
.save i(xdut.x1.v_isnk)
.save v(xdut.x1.Vpre)
.save i(xdut.x1.v_iPreCharge)
.save v(clk)
.save v(reset)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

unset askquit

optran 0 0 0 1n 1u 0

tran 100n 3u
write
quit


.endc

.end
