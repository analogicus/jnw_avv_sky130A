*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_bandgap_lpe.spi
#else
.include ../../../work/xsch/TB_bandgap.spice
#endif



*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option GMIN=1e-13 TNOM=25 
.option TEMP=20

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param PERIOD_CLK = {50e-9}
.param PW_CLK = PERIOD_CLK/2
.param T_START = PERIOD_CLK*4
.param T_RESET = {T_START + PERIOD_CLK + PW_CLK}
.param T_RESET_F = {T_RESET + 1n}
.param nbpt = 9*(8+5+2)

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS    0   dc 0
VDD  vdd    0   dc {AVDD}
VRST reset  0   dc 0
VCLK clk    0   dc 0 pulse (0 {AVDD} {T_START} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(clk)
.save v(vdd)
.save v(vss)
.save v(pa)
.save v(pb)
.save v(pc)
.save v(pd)
.save v(pi1)
.save v(pi2)
.save v(pii1)
.save v(pii2)
.save v(vref)
.save v(snk)
.save v(src)
.save v(xdut.vctrl)
.save v(xdut.pbias)
.save v(xdut.nbias)
.save v(xdut.vp)
.save v(xdut.vn)
.save v(reset)
.save v(cmp)
* .save v(valid)
* .save v(rst)
.save v(xdut.x3.snk_gate)
.save v(xdut.x3.src_gate_n)
.save v(xdut.x3.src_cap)
.save v(xdut.x3.snk_cap)
* .save v(xdut.x3.Vpre)
* .save i(xdut.v_nbias)
* .save i(xdut.v_pbias)
.save i(xdut.x2.vipmos)
.save v(xdut.x2.Hcharge)
.save v(xdut.x2.Lcharge)
.save v(xdut.x2.outRes)
.save v(xdut.x2.BD)
.save v(xdut.x2.SD)
.save v(xdut.x2.SDM)
.save v(xdut.x2.BDM)
.save v(xdut.x2.VbeSD)
.save v(xdut.x2.VbeBD)
.save v(xdut.x2.vpm)
.save v(xdut.x2.vnm)
.save i(vdd)
.save i(vss)
.save v(xdut.x1.ip)
.save v(xdut.x1.in)
.save v(xdut.x1.VipDrain)
.save v(xdut.x1.VinDrain)
.save v(xdut.x1.pre_vout)
.save v(xdut.x1.pre_voutn)
.save v(xdut.x1.vip)
.save v(xdut.x1.vin)
.save v(cmp_p1)
.save v(cmp_p2)


#ifdef debug
     .save all
     .option savecurrents
#endif

* .save all
* .option savecurrents


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

unset askquit

optran 0 0 0 100p 1.5u 0


set fend = .raw
* set debug = debug_


* tran 200n 40u


foreach vtemp 20
* foreach vtemp -40 -30 -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120 125
* foreach vtemp -40 -20 0 20 40 60 80 100 125
  option temp=$vtemp
  tran 1000n 40u
  write {cicname}_$vtemp$fend
end


write
quit


.endc

.end
