*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_bandgap_lpe.spi
#else
.include ../../../work/xsch/TB_bandgap.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

.param Vhigh = 1.8
.param Vlow = 0
.param low_th = 0.1
.param high_th = 1.7

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  vdd  VSS   dc 1.8

Vsrc  src  cmp   dc 0    
Vsnk  snk  cmp   dc 0   

*Vsrc  src  VSS   pulse 0 1.8 0 2n 2n 5u 10u 3 
*Vsnk  snk  VSS   pulse 0 1.8 0 2n 2n 5u 10u 3

VPA   PA   VSS   dc 0          
VPB   PB   VSS   dc 0          
VPC   PC   VSS   dc 0          
VPD   PD   VSS   dc 0          

* Pulse train and single pulse:
*VPI1  PI1  VSS   pulse 0 1.8 0 2n 2n 50u 100u 5           
*VPI1  PI1  VSS   pulse 0 1.8 100u 2n 2n 50u 100u 1

*VPI1  PI1  VSS   dc 1.8           
*VPI2  PI2  VSS   dc 1.8           

BPI1  PI1  VSS   V = V(cmp) < {low_th} ? {Vlow} :
    + V(cmp) > {high_th} ? {Vhigh}
BPI2  PI2  VSS   V = V(cmp) < {low_th} ? {Vlow} :
    + V(cmp) > {high_th} ? {Vhigh} : V(cmp)


VPII1 PII1 VSS   dc 0
VPII2 PII2 PII1  dc 0             

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1000n 30u
write
quit


.endc

.end
