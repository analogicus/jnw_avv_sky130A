*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CMP_lpe.spi
#else
.include ../../../work/xsch/CMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS     VSS   0     dc 0
VDD     VDD   VSS   dc 3
Vip     Vip   VSS   pwl 0 1.48 2 1.52
*Vip     Vip   VSS   dc 0
Vin     vin   VSS   dc 1.5
Itail   VDD   itail dc 12.5u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

tran 5m 2
*dc Vip 1.48 1.52 0.0001
write 
quit


.endc

.end
