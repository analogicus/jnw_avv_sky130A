*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_CMP_lpe.spi
#else
.include ../../../work/xsch/TB_CMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {1.8}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS  pwl 0 0 10n {AVDD}
Vip  vip   VSS   pwl 0 0.89 1000m 0.91 2000m 0.89 3000m 0.91 4000m 0.89
Vin  vin   VSS   pwl 0 0.91 1000m 0.89 2000m 0.91 3000m 0.89 4000m 0.91

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(cmp)
.save v(vip)
.save v(vin)
.save v(VDD)
.save v(VSS)
.save v(pbias)
.save v(nbias)



*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1m 4000m
write
quit


.endc

.end
