*Automatic generated instance fron ../../tech/scripts/gensvinst tmpDig
adut [clk
+ reset
+ cmp
+ ]
+ [PI1
+ PI2
+ PII1
+ dummy
+ PII2
+ PA
+ PB
+ PC
+ PD
+ s_BG2CMP
+ s_BgCtrl
+ s_PtatCtrl
+ s_Cap2CMP
+ s_Ref2CMP
+ s_CapRst
+ s_PtatOut
+ s_Rdiscon_N
+ src_n
+ snk
+ cmp_p1
+ cmp_p2
+ rst
+ valid
+ preChrg
+ setupBias
+ ] null dut
.model dut d_cosim simulation="../tmpDig.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 reset 0 1G
Rsvi2 cmp 0 1G

* Outputs
Rsvi3 PI1 0 1G
Rsvi4 PI2 0 1G
Rsvi5 PII1 0 1G
Rsvi6 dummy 0 1G
Rsvi7 PII2 0 1G
Rsvi8 PA 0 1G
Rsvi9 PB 0 1G
Rsvi10 PC 0 1G
Rsvi11 PD 0 1G
Rsvi12 s_BG2CMP 0 1G
Rsvi13 s_BgCtrl 0 1G
Rsvi14 s_PtatCtrl 0 1G
Rsvi15 s_Cap2CMP 0 1G
Rsvi16 s_Ref2CMP 0 1G
Rsvi17 s_CapRst 0 1G
Rsvi18 s_PtatOut 0 1G
Rsvi19 s_Rdiscon_N 0 1G
Rsvi20 src_n 0 1G
Rsvi21 snk 0 1G
Rsvi22 cmp_p1 0 1G
Rsvi23 cmp_p2 0 1G
Rsvi24 rst 0 1G
Rsvi25 valid 0 1G
Rsvi26 preChrg 0 1G
Rsvi27 setupBias 0 1G

.save v(PI1)

.save v(PI2)

.save v(PII1)

.save v(dummy)

.save v(PII2)

.save v(PA)

.save v(PB)

.save v(PC)

.save v(PD)

.save v(s_BG2CMP)

.save v(s_BgCtrl)

.save v(s_PtatCtrl)

.save v(s_Cap2CMP)

.save v(s_Ref2CMP)

.save v(s_CapRst)

.save v(s_PtatOut)

.save v(s_Rdiscon_N)

.save v(src_n)

.save v(snk)

.save v(cmp_p1)

.save v(cmp_p2)

.save v(rst)

.save v(valid)

.save v(preChrg)

.save v(setupBias)

