*Automatic generated instance fron ../../tech/scripts/genxdut tmpDig
adut [clk
+ reset
+ cmp
+ ]
+ [PI1
+ PI2
+ PII1
+ dummy
+ PII2
+ PA
+ PB
+ PC
+ PD
+ src_n
+ snk
+ cmp_p1
+ cmp_p2
+ sample
+ rst
+ valid
+ preChrg
+ setupBias
+ ] null dut
.model dut d_cosim simulation="../tmpDig.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 reset 0 1G
Rsvi2 cmp 0 1G

* Outputs
Rsvi3 PI1 0 1G
Rsvi4 PI2 0 1G
Rsvi5 PII1 0 1G
Rsvi6 dummy 0 1G
Rsvi7 PII2 0 1G
Rsvi8 PA 0 1G
Rsvi9 PB 0 1G
Rsvi10 PC 0 1G
Rsvi11 PD 0 1G
Rsvi12 src_n 0 1G
Rsvi13 snk 0 1G
Rsvi14 cmp_p1 0 1G
Rsvi15 cmp_p2 0 1G
Rsvi16 sample 0 1G
Rsvi17 rst 0 1G
Rsvi18 valid 0 1G
Rsvi19 preChrg 0 1G
Rsvi20 setupBias 0 1G

.save v(PI1)

.save v(PI2)

.save v(PII1)

.save v(dummy)

.save v(PII2)

.save v(PA)

.save v(PB)

.save v(PC)

.save v(PD)

.save v(src_n)

.save v(snk)

.save v(cmp_p1)

.save v(cmp_p2)

.save v(sample)

.save v(rst)

.save v(valid)

.save v(preChrg)

.save v(setupBias)

