*Automatic generated instance fron ../../tech/scripts/genxdut tmpDig
adut [clk
+ reset
+ cmp
+ ]
+ [PI1
+ PI2
+ PII1
+ PII2
+ PA
+ PB
+ PC
+ PD
+ src
+ snk
+ rst
+ valid
+ ] null dut
.model dut d_cosim simulation="../tmpDig.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 reset 0 1G
Rsvi2 cmp 0 1G

* Outputs
Rsvi3 PI1 0 1G
Rsvi4 PI2 0 1G
Rsvi5 PII1 0 1G
Rsvi6 PII2 0 1G
Rsvi7 PA 0 1G
Rsvi8 PB 0 1G
Rsvi9 PC 0 1G
Rsvi10 PD 0 1G
Rsvi11 src 0 1G
Rsvi12 snk 0 1G
Rsvi13 rst 0 1G
Rsvi14 valid 0 1G

.save v(PI1)

.save v(PI2)

.save v(PII1)

.save v(PII2)

.save v(PA)

.save v(PB)

.save v(PC)

.save v(PD)

.save v(src)

.save v(snk)

.save v(rst)

.save v(valid)

