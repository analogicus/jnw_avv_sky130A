*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bgTest_lpe.spi
#else
.include ../../../work/xsch/bgTest.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=25 GMIN=1e-15 reltol=1e-3
.option TEMP=20

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc 1.8

VA  A  0  pulse(0 1.8 0 10p 10p 300n 600n)
VB  B  0  dc 0.63055

* VA  A  0  pwl 0 0 50n 0 51n 1.8 150n 1.8 151n 0
* VB  B  0  pwl 0 0 100n 0 101n 1.8 200n 1.8 201n 0



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(vdd)
.save v(vss)
.save i(xdut.v_itot)
.save i(xdut.v_ip1)
.save i(xdut.v_ip2)
.save i(xdut.v_in1)
.save i(xdut.v_in2)
.save v(vref)
.save v(vp)
.save v(vn)
.save v(xdut.vctrl)
.save v(VBE)
.save v(A)
.save v(B)
.save v(xdut.y)
.save v(xdut.clk1)
.save v(xdut.clk2)
.save v(xdut.VBP)
.save v(xdut.VCP)
.save v(xdut.nbias)
.save v(xdut.pbias)
.save v(xdut.VbeBD)
.save v(xdut.vp)
.save v(xdut.bd)
.save v(xdut.bdm)
.save v(xdut.vpm)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


*dc TEMP -40 125 1
set fend = .raw


* foreach vtemp -40 -39 -38 -37 -36 -34 -32 -30 -28 -26 -24 -22 -20 -18 -16 -14 -12 -10 -8 -6
*   option temp=$vtemp
*   tran 10n 500n
*   write {cicname}_$vtemp$fend
* end

tran 0.5n 3u

write
quit


.endc

.end
