*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_leakage_lpe.spi
#else
.include ../../../work/xsch/TB_leakage.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  vss  0     dc 0
VDD  vdd  vss     dc {AVDD}

.ic v(xdut.x1.vn) = 0.6
.ic v(xdut.x1.vp) = 0.6
.ic v(xdut.x1.vref) = 0.6

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .save all
.save v(xdut.x1.vn)
.save v(xdut.x1.vp)
.save v(xdut.x1.vref)



*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1u 1m 0


tran 1n 10n 1p
write
quit


.endc

.end
