*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_charge_pump_lpe.spi
#else
.include ../../../work/xsch/TB_charge_pump.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  vdd  VSS   dc 1.8

Vsrc  src_n  VSS   pulse 0 1.8 0 2n 2n 50n 100n 7
Vsnk  snk  VSS   pulse 0 1.8 0 2n 2n 50n 100n 7
VpreChrg preChrg VSS dc 0

*Vsrc  src  VSS dc 0
*Vsnk  snk  VSS dc 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(vdd) 
.save v(vss)
.save v(src_n)
.save v(snk)
.save v(vctrl)
.save v(xdut.pbias)
.save v(xdut.nbias)
.save v(preChrg)
.save v(xdut.x1.snk_gate)
.save v(xdut.x1.src_n_gate)
.save v(xdut.x1.and_input)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

tran 2n 2u
write
quit


.endc

.end
