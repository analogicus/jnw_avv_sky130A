*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/bgTest_lpe.spi
#else
.include ../../../work/xsch/bgTest.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=25 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc 1.8



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(vdd)
.save v(vss)
.save i(xdut.v_itot)
.save i(xdut.v_ip1)
.save i(xdut.v_ip2)
.save i(xdut.v_in1)
.save i(xdut.v_in2)
.save v(vref)
.save v(vp)
.save v(vn)
.save v(xdut.vctrl)
.save v(VBE)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


*dc TEMP -40 125 1
tran 10n 10u
write
quit


.endc

.end
