*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CMP_lpe.spi
#else
.include ../../../work/xsch/CMP_v2.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS     VSS   0     dc 0
VDD     VDD   VSS   dc 1.8
*Vip     Vip   VSS   dc 0
Vip     vip   VSS   pwl 0 0.89 1000m 0.91 2000m 0.89
Vin     vin   VSS   pwl 0 0.91 1000m 0.89 2000m 0.91
*Vin     vin   VSS   dc 0.9
Itail   itail VSS   dc 12.5u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

tran 1m 2000m
*dc Vip 1.49 1.51 0.001
write 
quit


.endc

.end
