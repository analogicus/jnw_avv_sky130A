*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_bandgap_lpe.spi
#else
.include ../../../work/xsch/TB_bandgap.spice
#endif



*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option GMIN=1e-12 TNOM=25 reltol=1e-2
.option TEMP=20

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param PERIOD_CLK = {50e-9}
.param PW_CLK = PERIOD_CLK/2
.param T_START = PERIOD_CLK*4
.param T_RESET = {T_START + PERIOD_CLK + PW_CLK}
.param T_RESET_F = {T_RESET + 1n}
.param nbpt = 9*(8+5+2)



*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS    0   dc 0
VDD  vdd    0   dc {AVDD}
VRST reset  0   pwl 0 0 25n 0 25.1n 1.8 75n 1.8 75.1n 0
VCLK clk    0   dc 0 pulse (0 {AVDD} {T_START} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
* VCLK clk    0   dc 0 pulse (0 {AVDD} {18.8m} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi
* .include ../output_tran/ic/tran_schgtkttttvt_20.txt

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(clk)
.save v(vdd)
.save v(vss)
.save v(pa)
.save v(pb)
.save v(pc)
.save v(pd)
.save v(pi1)
.save v(pi2)
.save v(pii1)
.save v(pii2)
.save v(vref)
.save v(s_BG2CMP)
.save v(s_BgCtrl)
.save v(s_PtatCtrl)
.save v(s_Cap2CMP)
.save v(s_Ref2CMP)
.save v(s_CapRst)
.save v(s_PtatOut)
.save v(s_Rdiscon_N)
.save v(snk)
.save v(src_n)
.save v(xdut.vctrl)
.save v(xdut.pbias)
.save v(xdut.nbias)
.save v(xdut.vp)
.save v(xdut.vn)
.save i(xdut.x7.vIptat)
.save v(reset)
.save v(cmp)
.save v(tmpPulse)
* .save v(valid)
* .save v(rst)
.save v(xdut.x3.snk_gate)
.save v(xdut.x3.src_gate_n)
.save v(xdut.x3.src_cap)
.save v(xdut.x3.snk_cap)
.save v(xdut.x3.Vpre)
.save v(xdut.x3.vPtatCtrl)
.save v(xdut.x3.vBgCtrl)
* .save i(xdut.v_nbias)
* .save i(xdut.v_pbias)
.save i(xdut.x2.vipmos)
.save v(xdut.x2.Hcharge)
.save v(xdut.x2.Lcharge)
.save v(xdut.x2.vref)
.save v(xdut.x2.outRes)
.save v(xdut.x2.vpm)
.save v(xdut.x2.vnm)
.save v(xdut.x2.pmosDrain)
.save v(xdut.x2.cascDrain)
.save v(xdut.x2.pcasc)
.save v(xdut.OTAout)
.save v(xdut.OTAvip)
.save i(vdd)
.save i(vss)
.save v(xdut.x1.ip)
.save v(xdut.x1.in)
.save v(xdut.x1.VipDrain)
.save v(xdut.x1.VinDrain)
.save v(xdut.x1.inSource)
.save v(xdut.x1.pre_vout)
.save v(xdut.x1.pre_voutn)
.save v(xdut.x1.vip)
.save v(xdut.x1.vin)
.save v(xdut.x1.inShifted)
.save v(xdut.x1.ipShifted)
.save v(xdut.x1.in_intermediate)
.save v(xdut.x1.ip_intermediate)
.save i(xdut.x1.vibigdiode)
.save v(cmp_p1)
.save v(cmp_p2)
.save v(xdut.Vcap)
.save v(xdut.vin)
.save v(xdut.vip)
.save v(xdut.x7.Vcap2)
.save v(xdut.x7.Vcap1)
.save v(xdut.x7.rstCap1)
.save v(xdut.x7.rstCap2)
.save v(tmpCountRst_out)
.save v(tmpcount_out1)
.save v(tmpcount_out2)
.save v(tmpCount_out3)
.save v(tmpCount_out4)
.save v(count_out)
.save v(tmpSampleCount_out)

#ifdef debug
     .save all
     .option savecurrents
#endif

* .save all
* .option savecurrents


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

unset askquit

optran 0 0 0 100p 1.5u 0


set fend = .raw
set icend = .txt


******* Tempsens simulation ***********
foreach vtemp 20
* foreach vtemp -40 0 40 80 125
* foreach vtemp -40 20 0 -20 40 60 80 100 125
  option temp=$vtemp
  tran 1n 120u
*   wrnodev ic/{cicname}_$vtemp$icend
  write {cicname}_$vtemp$fend
end
****************************************



* *********** Leakage simulation ***********
* foreach vtemp 20
*   option temp=$vtemp
*   tran 1000n 18.91m
*   write {cicname}_$vtemp$fend
* end
* *******************************************




write
quit


.endc
.end
